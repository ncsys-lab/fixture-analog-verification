.lib "/home/will/Desktop/AchourLab/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice" tt


.subckt LDO_COMPARATOR_LATCH vgnd vpwr VREF VREG CLK outp outn
R0 vnb vgnd 0
R1 vpb vpwr 0
R2 a_512_1261# outp 0
R3 a_519_81# outn 0
X0 a_612_1321# a_512_1261# a_123_187# vnb sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u nf=5
X1 a_612_1321# VREF a_519_81# vnb sky130_fd_pr__nfet_g5v0d10v5 w=10e+06u l=500000u nf=10
X2 vpwr OUT a_3401_885# vpb sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_519_81# a_512_1261# vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 w=10e+06u l=500000u 
X4 a_512_1261# a_519_81# vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 w=10e+06u l=500000u 
X5 a_519_81# CLK vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u 
X6 vpwr CLK a_512_1261# vpb sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u 
X7 a_619_107# VREG a_512_1261# vnb sky130_fd_pr__nfet_g5v0d10v5 w=10e+06u l=500000u
X8 OUT a_512_1261# vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_123_187# a_519_81# a_619_107# vnb sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u 
X10 a_3401_111# a_512_1261# vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 OUT a_3401_885# a_3401_111# vnb sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 a_3401_1367# a_519_81# vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 a_3401_885# a_519_81# vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_3401_885# OUT a_3401_1367# vnb sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 vgnd CLK a_123_187# vnb sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 vpwr a_3401_885# OUT vpb sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends
