* Automatically generated file.
.include /home/will/Desktop/AchourLab/fixture-analog-verification/tests/spice/LDO_COMPARATOR_LATCH.spice
X0 vgnd vpwr vref vreg clk outp outn LDO_COMPARATOR_LATCH
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __vpwr_v vpwr __vpwr_s 0 inout_sw_mod
V2 __vpwr_v 0 DC 3.3 PWL(0 3.3 0.00015026400000000008 3.3)
V3 __vpwr_s 0 DC 1 PWL(0 1 0.00015026400000000008 1)
X4 __vgnd_v vgnd __vgnd_s 0 inout_sw_mod
V5 __vgnd_v 0 DC 0 PWL(0 0 0.00015026400000000008 0)
V6 __vgnd_s 0 DC 1 PWL(0 1 0.00015026400000000008 1)
X7 __CLK_v CLK __CLK_s 0 inout_sw_mod
V8 __CLK_v 0 DC 0 PWL(0 0 4.9999999999999996e-06 0 5.000199999999999e-06 3.3 5.008799999999999e-06 3.3 5.008999999999999e-06 0 1.0008799999999998e-05 0 1.0008999999999999e-05 3.3 1.0017599999999999e-05 3.3 1.00178e-05 0 1.5017599999999998e-05 0 1.5017799999999999e-05 3.3 1.5026399999999999e-05 3.3 1.50266e-05 0 2.00264e-05 0 2.00266e-05 3.3 2.0035199999999998e-05 3.3 2.0035399999999998e-05 0 2.5035199999999997e-05 0 2.5035399999999998e-05 3.3 2.5043999999999996e-05 3.3 2.5044199999999996e-05 0 3.0043999999999996e-05 0 3.0044199999999996e-05 3.3 3.0052799999999995e-05 3.3 3.0052999999999995e-05 0 3.50528e-05 0 3.5053e-05 3.3 3.5061599999999996e-05 3.3 3.50618e-05 0 4.0061599999999996e-05 0 4.0061799999999996e-05 3.3 4.0070399999999995e-05 3.3 4.0070599999999995e-05 0 4.5070399999999995e-05 0 4.5070599999999995e-05 3.3 4.5079199999999994e-05 3.3 4.5079399999999994e-05 0 5.007919999999999e-05 0 5.0079399999999994e-05 3.3 5.008799999999999e-05 3.3 5.008819999999999e-05 0 5.508799999999999e-05 0 5.508819999999999e-05 3.3 5.509679999999999e-05 3.3 5.509699999999999e-05 0 6.009679999999999e-05 0 6.009699999999999e-05 3.3 6.010559999999999e-05 3.3 6.010579999999999e-05 0 6.51056e-05 0 6.51058e-05 3.3 6.51144e-05 3.3 6.51146e-05 0 7.01144e-05 0 7.01146e-05 3.3 7.01232e-05 3.3 7.012340000000001e-05 0 7.51232e-05 0 7.51234e-05 3.3 7.513200000000001e-05 3.3 7.513220000000001e-05 0 8.013200000000001e-05 0 8.013220000000001e-05 3.3 8.014080000000002e-05 3.3 8.014100000000002e-05 0 8.514080000000002e-05 0 8.514100000000002e-05 3.3 8.514960000000002e-05 3.3 8.514980000000002e-05 0 9.014960000000002e-05 0 9.014980000000002e-05 3.3 9.015840000000003e-05 3.3 9.015860000000003e-05 0 9.515840000000003e-05 0 9.515860000000003e-05 3.3 9.516720000000003e-05 3.3 9.516740000000003e-05 0 0.00010016720000000003 0 0.00010016740000000003 3.3 0.00010017600000000004 3.3 0.00010017620000000004 0 0.00010517600000000004 0 0.00010517620000000004 3.3 0.00010518480000000004 3.3 0.00010518500000000004 0 0.00011018480000000004 0 0.00011018500000000004 3.3 0.00011019360000000005 3.3 0.00011019380000000005 0 0.00011519360000000005 0 0.00011519380000000005 3.3 0.00011520240000000005 3.3 0.00011520260000000005 0 0.00012020240000000005 0 0.00012020260000000005 3.3 0.00012021120000000006 3.3 0.00012021140000000006 0 0.00012521120000000006 0 0.00012521140000000005 3.3 0.00012522000000000005 3.3 0.00012522020000000004 0 0.00013022000000000006 0 0.00013022020000000005 3.3 0.00013022880000000006 3.3 0.00013022900000000004 0 0.00013522880000000007 0 0.00013522900000000006 3.3 0.00013523760000000006 3.3 0.00013523780000000005 0 0.00014023760000000008 0 0.00014023780000000006 3.3 0.00014024640000000007 3.3 0.00014024660000000005 0 0.00014524640000000008 0 0.00014524660000000007 3.3 0.00014525520000000007 3.3 0.00014525540000000006 0 0.00015025520000000009 0 0.00015025540000000007 3.3 0.00015026400000000008 3.3)
V9 __CLK_s 0 DC 1 PWL(0 1 4.9999999999999996e-06 1 5.000199999999999e-06 1 5.008799999999999e-06 1 5.008999999999999e-06 1 1.0008799999999998e-05 1 1.0008999999999999e-05 1 1.0017599999999999e-05 1 1.00178e-05 1 1.5017599999999998e-05 1 1.5017799999999999e-05 1 1.5026399999999999e-05 1 1.50266e-05 1 2.00264e-05 1 2.00266e-05 1 2.0035199999999998e-05 1 2.0035399999999998e-05 1 2.5035199999999997e-05 1 2.5035399999999998e-05 1 2.5043999999999996e-05 1 2.5044199999999996e-05 1 3.0043999999999996e-05 1 3.0044199999999996e-05 1 3.0052799999999995e-05 1 3.0052999999999995e-05 1 3.50528e-05 1 3.5053e-05 1 3.5061599999999996e-05 1 3.50618e-05 1 4.0061599999999996e-05 1 4.0061799999999996e-05 1 4.0070399999999995e-05 1 4.0070599999999995e-05 1 4.5070399999999995e-05 1 4.5070599999999995e-05 1 4.5079199999999994e-05 1 4.5079399999999994e-05 1 5.007919999999999e-05 1 5.0079399999999994e-05 1 5.008799999999999e-05 1 5.008819999999999e-05 1 5.508799999999999e-05 1 5.508819999999999e-05 1 5.509679999999999e-05 1 5.509699999999999e-05 1 6.009679999999999e-05 1 6.009699999999999e-05 1 6.010559999999999e-05 1 6.010579999999999e-05 1 6.51056e-05 1 6.51058e-05 1 6.51144e-05 1 6.51146e-05 1 7.01144e-05 1 7.01146e-05 1 7.01232e-05 1 7.012340000000001e-05 1 7.51232e-05 1 7.51234e-05 1 7.513200000000001e-05 1 7.513220000000001e-05 1 8.013200000000001e-05 1 8.013220000000001e-05 1 8.014080000000002e-05 1 8.014100000000002e-05 1 8.514080000000002e-05 1 8.514100000000002e-05 1 8.514960000000002e-05 1 8.514980000000002e-05 1 9.014960000000002e-05 1 9.014980000000002e-05 1 9.015840000000003e-05 1 9.015860000000003e-05 1 9.515840000000003e-05 1 9.515860000000003e-05 1 9.516720000000003e-05 1 9.516740000000003e-05 1 0.00010016720000000003 1 0.00010016740000000003 1 0.00010017600000000004 1 0.00010017620000000004 1 0.00010517600000000004 1 0.00010517620000000004 1 0.00010518480000000004 1 0.00010518500000000004 1 0.00011018480000000004 1 0.00011018500000000004 1 0.00011019360000000005 1 0.00011019380000000005 1 0.00011519360000000005 1 0.00011519380000000005 1 0.00011520240000000005 1 0.00011520260000000005 1 0.00012020240000000005 1 0.00012020260000000005 1 0.00012021120000000006 1 0.00012021140000000006 1 0.00012521120000000006 1 0.00012521140000000005 1 0.00012522000000000005 1 0.00012522020000000004 1 0.00013022000000000006 1 0.00013022020000000005 1 0.00013022880000000006 1 0.00013022900000000004 1 0.00013522880000000007 1 0.00013522900000000006 1 0.00013523760000000006 1 0.00013523780000000005 1 0.00014023760000000008 1 0.00014023780000000006 1 0.00014024640000000007 1 0.00014024660000000005 1 0.00014524640000000008 1 0.00014524660000000007 1 0.00014525520000000007 1 0.00014525540000000006 1 0.00015025520000000009 1 0.00015025540000000007 1 0.00015026400000000008 1)
X10 __VREG_v VREG __VREG_s 0 inout_sw_mod
V11 __VREG_v 0 DC 0 PWL(0 0 2.4999999999999998e-06 0 2.5002e-06 2.9047209617947485 7.508799999999999e-06 2.9047209617947485 7.508999999999999e-06 2.909934304043511 1.2517599999999999e-05 2.909934304043511 1.2517799999999999e-05 2.9008868679423943 1.75264e-05 2.9008868679423943 1.75266e-05 2.919179550430877 2.2535199999999997e-05 2.919179550430877 2.2535399999999998e-05 2.915101084016703 2.7543999999999996e-05 2.915101084016703 2.7544199999999996e-05 2.9307336001634963 3.25528e-05 2.9307336001634963 3.2553e-05 2.922877742154756 3.7561599999999996e-05 2.922877742154756 3.75618e-05 2.9261920057677187 4.2570399999999995e-05 2.9261920057677187 4.2570599999999995e-05 2.9382892004877843 4.757919999999999e-05 2.9382892004877843 4.7579399999999994e-05 2.93533631892362 5.258799999999999e-05 2.93533631892362 5.258819999999999e-05 2.946196999145991 5.759679999999999e-05 2.946196999145991 5.759699999999999e-05 2.955531578481312 6.260559999999999e-05 2.955531578481312 6.260579999999999e-05 2.958400676684816 6.76144e-05 2.958400676684816 6.76146e-05 2.9493918521705322 7.26232e-05 2.9493918521705322 7.26234e-05 2.9500396918380694 7.7632e-05 2.9500396918380694 7.76322e-05 2.9694717577517027 8.264080000000001e-05 2.9694717577517027 8.264100000000001e-05 2.9789098060649986 8.764960000000002e-05 2.9789098060649986 8.764980000000002e-05 2.9706351849278274 9.265840000000002e-05 2.9706351849278274 9.265860000000002e-05 2.9757553695608134 9.766720000000003e-05 2.9757553695608134 9.766740000000003e-05 2.9658821149325254 0.00010267600000000003 2.9658821149325254 0.00010267620000000003 2.990167447506655 0.00010768480000000004 2.990167447506655 0.00010768500000000004 2.9899818745365 0.00011269360000000004 2.9899818745365 0.00011269380000000004 2.9821509414149547 0.00011770240000000005 2.9821509414149547 0.00011770260000000005 2.9981259231863464 0.00012271120000000005 2.9981259231863464 0.00012271140000000004 2.9836421466600234 0.00012772000000000006 2.9836421466600234 0.00012772020000000004 2.9284487393162646 0.00013272880000000006 2.9284487393162646 0.00013272900000000005 2.993985244981111 0.00013773760000000007 2.993985244981111 0.00013773780000000006 2.9409210161165324 0.00014274640000000007 2.9409210161165324 0.00014274660000000006 2.911861763278611 0.00014775520000000008 2.911861763278611 0.00014775540000000007 2.960762898134129 0.00015026400000000008 2.960762898134129)
V12 __VREG_s 0 DC 1 PWL(0 1 2.4999999999999998e-06 1 2.5002e-06 1 7.508799999999999e-06 1 7.508999999999999e-06 1 1.2517599999999999e-05 1 1.2517799999999999e-05 1 1.75264e-05 1 1.75266e-05 1 2.2535199999999997e-05 1 2.2535399999999998e-05 1 2.7543999999999996e-05 1 2.7544199999999996e-05 1 3.25528e-05 1 3.2553e-05 1 3.7561599999999996e-05 1 3.75618e-05 1 4.2570399999999995e-05 1 4.2570599999999995e-05 1 4.757919999999999e-05 1 4.7579399999999994e-05 1 5.258799999999999e-05 1 5.258819999999999e-05 1 5.759679999999999e-05 1 5.759699999999999e-05 1 6.260559999999999e-05 1 6.260579999999999e-05 1 6.76144e-05 1 6.76146e-05 1 7.26232e-05 1 7.26234e-05 1 7.7632e-05 1 7.76322e-05 1 8.264080000000001e-05 1 8.264100000000001e-05 1 8.764960000000002e-05 1 8.764980000000002e-05 1 9.265840000000002e-05 1 9.265860000000002e-05 1 9.766720000000003e-05 1 9.766740000000003e-05 1 0.00010267600000000003 1 0.00010267620000000003 1 0.00010768480000000004 1 0.00010768500000000004 1 0.00011269360000000004 1 0.00011269380000000004 1 0.00011770240000000005 1 0.00011770260000000005 1 0.00012271120000000005 1 0.00012271140000000004 1 0.00012772000000000006 1 0.00012772020000000004 1 0.00013272880000000006 1 0.00013272900000000005 1 0.00013773760000000007 1 0.00013773780000000006 1 0.00014274640000000007 1 0.00014274660000000006 1 0.00014775520000000008 1 0.00014775540000000007 1 0.00015026400000000008 1)
X13 __VREF_v VREF __VREF_s 0 inout_sw_mod
V14 __VREF_v 0 DC 0 PWL(0 0 2.4999999999999998e-06 0 2.5002e-06 1.5041266413692287 7.508799999999999e-06 1.5041266413692287 7.508999999999999e-06 1.5461988908320965 1.2517599999999999e-05 1.5461988908320965 1.2517799999999999e-05 1.5960636405794029 1.75264e-05 1.5960636405794029 1.75266e-05 1.6520180940598324 2.2535199999999997e-05 1.6520180940598324 2.2535399999999998e-05 1.6688771270276126 2.7543999999999996e-05 1.6688771270276126 2.7544199999999996e-05 1.5158894214480483 3.25528e-05 1.5158894214480483 3.2553e-05 1.5502061097477178 3.7561599999999996e-05 1.5502061097477178 3.75618e-05 1.617582521047602 4.2570399999999995e-05 1.617582521047602 4.2570599999999995e-05 1.6535550782234107 4.757919999999999e-05 1.6535550782234107 4.7579399999999994e-05 1.6664478539339747 5.258799999999999e-05 1.6664478539339747 5.258819999999999e-05 1.5300526827310168 5.759679999999999e-05 1.5300526827310168 5.759699999999999e-05 1.5761239562131026 6.260559999999999e-05 1.5761239562131026 6.260579999999999e-05 1.5823124867369311 6.76144e-05 1.5823124867369311 6.76146e-05 1.6379120388404393 7.26232e-05 1.6379120388404393 7.26234e-05 1.6780744046464209 7.7632e-05 1.6780744046464209 7.76322e-05 1.5084535908119745 8.264080000000001e-05 1.5084535908119745 8.264100000000001e-05 1.5706430167370349 8.764960000000002e-05 1.5706430167370349 8.764980000000002e-05 1.5926715814581331 9.265840000000002e-05 1.5926715814581331 9.265860000000002e-05 1.6314473360337178 9.766720000000003e-05 1.6314473360337178 9.766740000000003e-05 1.6969608817644726 0.00010267600000000003 1.6969608817644726 0.00010267620000000003 1.5255192805750897 0.00010768480000000004 1.5255192805750897 0.00010768500000000004 1.5590805735639108 0.00011269360000000004 1.5590805735639108 0.00011269380000000004 1.6040681546191031 0.00011770240000000005 1.6040681546191031 0.00011770260000000005 1.6205765129209633 0.00012271120000000005 1.6205765129209633 0.00012271140000000004 1.6883513432738653 0.00012772000000000006 1.6883513432738653 0.00012772020000000004 1.6089522884361478 0.00013272880000000006 1.6089522884361478 0.00013272900000000005 1.5613511374411493 0.00013773760000000007 1.5613511374411493 0.00013773780000000006 1.6449796178732696 0.00014274640000000007 1.6449796178732696 0.00014274660000000006 1.680673196258119 0.00014775520000000008 1.680673196258119 0.00014775540000000007 1.5374362138341913 0.00015026400000000008 1.5374362138341913)
V15 __VREF_s 0 DC 1 PWL(0 1 2.4999999999999998e-06 1 2.5002e-06 1 7.508799999999999e-06 1 7.508999999999999e-06 1 1.2517599999999999e-05 1 1.2517799999999999e-05 1 1.75264e-05 1 1.75266e-05 1 2.2535199999999997e-05 1 2.2535399999999998e-05 1 2.7543999999999996e-05 1 2.7544199999999996e-05 1 3.25528e-05 1 3.2553e-05 1 3.7561599999999996e-05 1 3.75618e-05 1 4.2570399999999995e-05 1 4.2570599999999995e-05 1 4.757919999999999e-05 1 4.7579399999999994e-05 1 5.258799999999999e-05 1 5.258819999999999e-05 1 5.759679999999999e-05 1 5.759699999999999e-05 1 6.260559999999999e-05 1 6.260579999999999e-05 1 6.76144e-05 1 6.76146e-05 1 7.26232e-05 1 7.26234e-05 1 7.7632e-05 1 7.76322e-05 1 8.264080000000001e-05 1 8.264100000000001e-05 1 8.764960000000002e-05 1 8.764980000000002e-05 1 9.265840000000002e-05 1 9.265860000000002e-05 1 9.766720000000003e-05 1 9.766740000000003e-05 1 0.00010267600000000003 1 0.00010267620000000003 1 0.00010768480000000004 1 0.00010768500000000004 1 0.00011269360000000004 1 0.00011269380000000004 1 0.00011770240000000005 1 0.00011770260000000005 1 0.00012271120000000005 1 0.00012271140000000004 1 0.00012772000000000006 1 0.00012772020000000004 1 0.00013272880000000006 1 0.00013272900000000005 1 0.00013773760000000007 1 0.00013773780000000006 1 0.00014274640000000007 1 0.00014274660000000006 1 0.00014775520000000008 1 0.00014775540000000007 1 0.00015026400000000008 1)
.tran 1e-10 0.00015026400000000008
.control
run
set filetype=binary
write
exit
.endc
.probe V(vpwr) V(outn) V(VREG) V(CLK) V(VREF) V(outp) V(vgnd)
.end
