* Automatically generated file.
.include /home/will/Desktop/AchourLab/fixture-analog-verification/tests/spice/LDO_COMPARATOR_LATCH.spice
X0 vgnd vpwr vref vreg clk outp outn LDO_COMPARATOR_LATCH
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __vpwr_v vpwr __vpwr_s 0 inout_sw_mod
V2 __vpwr_v 0 DC 3.3 PWL(0 3.3 0.00012199999999999978 3.3)
V3 __vpwr_s 0 DC 1 PWL(0 1 0.00012199999999999978 1)
X4 __vgnd_v vgnd __vgnd_s 0 inout_sw_mod
V5 __vgnd_v 0 DC 0 PWL(0 0 0.00012199999999999978 0)
V6 __vgnd_s 0 DC 1 PWL(0 1 0.00012199999999999978 1)
X7 __CLK_v CLK __CLK_s 0 inout_sw_mod
V8 __CLK_v 0 DC 0 PWL(0 0 9.999999999999999e-06 0 1.00002e-05 3.3 3.699999999999999e-05 3.3 3.700019999999999e-05 0 3.799999999999999e-05 0 3.800019999999999e-05 0 3.8999999999999986e-05 0 3.9000199999999986e-05 0 3.999999999999998e-05 0 4.000019999999998e-05 0 4.099999999999998e-05 0 4.100019999999998e-05 0 4.199999999999998e-05 0 4.200019999999998e-05 0 4.2999999999999975e-05 0 4.3000199999999975e-05 0 4.399999999999997e-05 0 4.400019999999997e-05 0 4.499999999999997e-05 0 4.500019999999997e-05 0 4.5999999999999966e-05 0 4.6000199999999967e-05 0 4.699999999999996e-05 0 4.7000199999999964e-05 3.3 4.799999999999996e-05 3.3 4.800019999999996e-05 3.3 4.899999999999996e-05 3.3 4.900019999999996e-05 3.3 4.9999999999999955e-05 3.3 5.0000199999999955e-05 3.3 5.099999999999995e-05 3.3 5.100019999999995e-05 3.3 5.199999999999995e-05 3.3 5.200019999999995e-05 3.3 5.2999999999999947e-05 3.3 5.300019999999995e-05 3.3 5.3999999999999944e-05 3.3 5.4000199999999944e-05 3.3 5.499999999999994e-05 3.3 5.500019999999994e-05 3.3 5.599999999999994e-05 3.3 5.600019999999994e-05 3.3 5.6999999999999935e-05 3.3 5.7000199999999936e-05 3.3 5.799999999999993e-05 3.3 5.800019999999993e-05 3.3 5.899999999999993e-05 3.3 5.900019999999993e-05 3.3 5.999999999999993e-05 3.3 6.000019999999993e-05 3.3 6.0999999999999924e-05 3.3 6.1000199999999925e-05 0 7.099999999999992e-05 0 7.100019999999992e-05 3.3 9.799999999999985e-05 3.3 9.800019999999985e-05 0 9.899999999999984e-05 0 9.900019999999985e-05 0 9.999999999999984e-05 0 0.00010000019999999984 0 0.00010099999999999984 0 0.00010100019999999984 0 0.00010199999999999984 0 0.00010200019999999984 0 0.00010299999999999983 0 0.00010300019999999983 0 0.00010399999999999983 0 0.00010400019999999983 0 0.00010499999999999983 0 0.00010500019999999983 0 0.00010599999999999983 0 0.00010600019999999983 0 0.00010699999999999982 0 0.00010700019999999982 0 0.00010799999999999982 0 0.00010800019999999982 3.3 0.00010899999999999982 3.3 0.00010900019999999982 3.3 0.00010999999999999981 3.3 0.00011000019999999981 3.3 0.00011099999999999981 3.3 0.00011100019999999981 3.3 0.00011199999999999981 3.3 0.00011200019999999981 3.3 0.0001129999999999998 3.3 0.0001130001999999998 3.3 0.0001139999999999998 3.3 0.0001140001999999998 3.3 0.0001149999999999998 3.3 0.0001150001999999998 3.3 0.0001159999999999998 3.3 0.0001160001999999998 3.3 0.0001169999999999998 3.3 0.0001170001999999998 3.3 0.00011799999999999979 3.3 0.00011800019999999979 3.3 0.00011899999999999979 3.3 0.00011900019999999979 3.3 0.00011999999999999979 3.3 0.00012000019999999979 3.3 0.00012099999999999978 3.3 0.00012100019999999978 3.3 0.00012199999999999978 3.3)
V9 __CLK_s 0 DC 1 PWL(0 1 9.999999999999999e-06 1 1.00002e-05 1 3.699999999999999e-05 1 3.700019999999999e-05 1 3.799999999999999e-05 1 3.800019999999999e-05 1 3.8999999999999986e-05 1 3.9000199999999986e-05 1 3.999999999999998e-05 1 4.000019999999998e-05 1 4.099999999999998e-05 1 4.100019999999998e-05 1 4.199999999999998e-05 1 4.200019999999998e-05 1 4.2999999999999975e-05 1 4.3000199999999975e-05 1 4.399999999999997e-05 1 4.400019999999997e-05 1 4.499999999999997e-05 1 4.500019999999997e-05 1 4.5999999999999966e-05 1 4.6000199999999967e-05 1 4.699999999999996e-05 1 4.7000199999999964e-05 1 4.799999999999996e-05 1 4.800019999999996e-05 1 4.899999999999996e-05 1 4.900019999999996e-05 1 4.9999999999999955e-05 1 5.0000199999999955e-05 1 5.099999999999995e-05 1 5.100019999999995e-05 1 5.199999999999995e-05 1 5.200019999999995e-05 1 5.2999999999999947e-05 1 5.300019999999995e-05 1 5.3999999999999944e-05 1 5.4000199999999944e-05 1 5.499999999999994e-05 1 5.500019999999994e-05 1 5.599999999999994e-05 1 5.600019999999994e-05 1 5.6999999999999935e-05 1 5.7000199999999936e-05 1 5.799999999999993e-05 1 5.800019999999993e-05 1 5.899999999999993e-05 1 5.900019999999993e-05 1 5.999999999999993e-05 1 6.000019999999993e-05 1 6.0999999999999924e-05 1 6.1000199999999925e-05 1 7.099999999999992e-05 1 7.100019999999992e-05 1 9.799999999999985e-05 1 9.800019999999985e-05 1 9.899999999999984e-05 1 9.900019999999985e-05 1 9.999999999999984e-05 1 0.00010000019999999984 1 0.00010099999999999984 1 0.00010100019999999984 1 0.00010199999999999984 1 0.00010200019999999984 1 0.00010299999999999983 1 0.00010300019999999983 1 0.00010399999999999983 1 0.00010400019999999983 1 0.00010499999999999983 1 0.00010500019999999983 1 0.00010599999999999983 1 0.00010600019999999983 1 0.00010699999999999982 1 0.00010700019999999982 1 0.00010799999999999982 1 0.00010800019999999982 1 0.00010899999999999982 1 0.00010900019999999982 1 0.00010999999999999981 1 0.00011000019999999981 1 0.00011099999999999981 1 0.00011100019999999981 1 0.00011199999999999981 1 0.00011200019999999981 1 0.0001129999999999998 1 0.0001130001999999998 1 0.0001139999999999998 1 0.0001140001999999998 1 0.0001149999999999998 1 0.0001150001999999998 1 0.0001159999999999998 1 0.0001160001999999998 1 0.0001169999999999998 1 0.0001170001999999998 1 0.00011799999999999979 1 0.00011800019999999979 1 0.00011899999999999979 1 0.00011900019999999979 1 0.00011999999999999979 1 0.00012000019999999979 1 0.00012099999999999978 1 0.00012100019999999978 1 0.00012199999999999978 1)
X10 __VREG_v VREG __VREG_s 0 inout_sw_mod
V11 __VREG_v 0 DC 0 PWL(0 0 1.1e-05 0 1.10002e-05 0.0 1.2e-05 0.0 1.20002e-05 0.0673469387755102 1.3000000000000001e-05 0.0673469387755102 1.3000200000000001e-05 0.1346938775510204 1.4000000000000001e-05 0.1346938775510204 1.4000200000000002e-05 0.20204081632653062 1.5000000000000002e-05 0.20204081632653062 1.5000200000000003e-05 0.2693877551020408 1.6000000000000003e-05 0.2693877551020408 1.6000200000000003e-05 0.33673469387755106 1.7000000000000003e-05 0.33673469387755106 1.7000200000000004e-05 0.40408163265306124 1.8000000000000004e-05 0.40408163265306124 1.8000200000000004e-05 0.4714285714285714 1.9000000000000004e-05 0.4714285714285714 1.9000200000000005e-05 0.5387755102040817 2.0000000000000005e-05 0.5387755102040817 2.0000200000000005e-05 0.6061224489795919 2.1000000000000006e-05 0.6061224489795919 2.1000200000000006e-05 0.6734693877551021 2.2000000000000006e-05 0.6734693877551021 2.2000200000000007e-05 0.7408163265306122 2.3000000000000007e-05 0.7408163265306122 2.3000200000000007e-05 0.8081632653061225 2.4000000000000007e-05 0.8081632653061225 2.4000200000000008e-05 0.8755102040816327 2.5000000000000008e-05 0.8755102040816327 2.500020000000001e-05 0.9428571428571428 2.600000000000001e-05 0.9428571428571428 2.600020000000001e-05 1.0102040816326532 2.700000000000001e-05 1.0102040816326532 2.700020000000001e-05 1.0775510204081633 2.800000000000001e-05 1.0775510204081633 2.800020000000001e-05 1.1448979591836734 2.900000000000001e-05 1.1448979591836734 2.900020000000001e-05 1.2122448979591838 3.000000000000001e-05 1.2122448979591838 3.000020000000001e-05 1.279591836734694 3.100000000000001e-05 1.279591836734694 3.100020000000001e-05 1.3469387755102042 3.2000000000000005e-05 1.3469387755102042 3.2000200000000006e-05 1.4142857142857144 3.3e-05 1.4142857142857144 3.30002e-05 1.4816326530612245 3.4e-05 1.4816326530612245 3.40002e-05 1.5489795918367348 3.5e-05 1.5489795918367348 3.50002e-05 1.616326530612245 3.5999999999999994e-05 1.616326530612245 3.6000199999999995e-05 1.683673469387755 3.699999999999999e-05 1.683673469387755 3.700019999999999e-05 1.7510204081632654 3.799999999999999e-05 1.7510204081632654 3.800019999999999e-05 1.8183673469387756 3.8999999999999986e-05 1.8183673469387756 3.9000199999999986e-05 1.8857142857142857 3.999999999999998e-05 1.8857142857142857 4.000019999999998e-05 1.953061224489796 4.099999999999998e-05 1.953061224489796 4.100019999999998e-05 2.0204081632653064 4.199999999999998e-05 2.0204081632653064 4.200019999999998e-05 2.0877551020408163 4.2999999999999975e-05 2.0877551020408163 4.3000199999999975e-05 2.1551020408163266 4.399999999999997e-05 2.1551020408163266 4.400019999999997e-05 2.222448979591837 4.499999999999997e-05 2.222448979591837 4.500019999999997e-05 2.289795918367347 4.5999999999999966e-05 2.289795918367347 4.6000199999999967e-05 2.357142857142857 4.699999999999996e-05 2.357142857142857 4.7000199999999964e-05 2.4244897959183676 4.799999999999996e-05 2.4244897959183676 4.800019999999996e-05 2.4918367346938775 4.899999999999996e-05 2.4918367346938775 4.900019999999996e-05 2.559183673469388 4.9999999999999955e-05 2.559183673469388 5.0000199999999955e-05 2.626530612244898 5.099999999999995e-05 2.626530612244898 5.100019999999995e-05 2.6938775510204085 5.199999999999995e-05 2.6938775510204085 5.200019999999995e-05 2.7612244897959184 5.2999999999999947e-05 2.7612244897959184 5.300019999999995e-05 2.8285714285714287 5.3999999999999944e-05 2.8285714285714287 5.4000199999999944e-05 2.895918367346939 5.499999999999994e-05 2.895918367346939 5.500019999999994e-05 2.963265306122449 5.599999999999994e-05 2.963265306122449 5.600019999999994e-05 3.0306122448979593 5.6999999999999935e-05 3.0306122448979593 5.7000199999999936e-05 3.0979591836734697 5.799999999999993e-05 3.0979591836734697 5.800019999999993e-05 3.1653061224489796 5.899999999999993e-05 3.1653061224489796 5.900019999999993e-05 3.23265306122449 5.999999999999993e-05 3.23265306122449 6.000019999999993e-05 3.3 6.0999999999999924e-05 3.3 6.1000199999999925e-05 0 7.199999999999992e-05 0 7.200019999999992e-05 0.0 7.299999999999992e-05 0.0 7.300019999999992e-05 0.0673469387755102 7.399999999999991e-05 0.0673469387755102 7.400019999999992e-05 0.1346938775510204 7.499999999999991e-05 0.1346938775510204 7.500019999999991e-05 0.20204081632653062 7.599999999999991e-05 0.20204081632653062 7.600019999999991e-05 0.2693877551020408 7.69999999999999e-05 0.2693877551020408 7.700019999999991e-05 0.33673469387755106 7.79999999999999e-05 0.33673469387755106 7.80001999999999e-05 0.40408163265306124 7.89999999999999e-05 0.40408163265306124 7.90001999999999e-05 0.4714285714285714 7.99999999999999e-05 0.4714285714285714 8.00001999999999e-05 0.5387755102040817 8.09999999999999e-05 0.5387755102040817 8.10001999999999e-05 0.6061224489795919 8.199999999999989e-05 0.6061224489795919 8.200019999999989e-05 0.6734693877551021 8.299999999999989e-05 0.6734693877551021 8.300019999999989e-05 0.7408163265306122 8.399999999999989e-05 0.7408163265306122 8.400019999999989e-05 0.8081632653061225 8.499999999999988e-05 0.8081632653061225 8.500019999999988e-05 0.8755102040816327 8.599999999999988e-05 0.8755102040816327 8.600019999999988e-05 0.9428571428571428 8.699999999999988e-05 0.9428571428571428 8.700019999999988e-05 1.0102040816326532 8.799999999999988e-05 1.0102040816326532 8.800019999999988e-05 1.0775510204081633 8.899999999999987e-05 1.0775510204081633 8.900019999999987e-05 1.1448979591836734 8.999999999999987e-05 1.1448979591836734 9.000019999999987e-05 1.2122448979591838 9.099999999999987e-05 1.2122448979591838 9.100019999999987e-05 1.279591836734694 9.199999999999986e-05 1.279591836734694 9.200019999999986e-05 1.3469387755102042 9.299999999999986e-05 1.3469387755102042 9.300019999999986e-05 1.4142857142857144 9.399999999999986e-05 1.4142857142857144 9.400019999999986e-05 1.4816326530612245 9.499999999999986e-05 1.4816326530612245 9.500019999999986e-05 1.5489795918367348 9.599999999999985e-05 1.5489795918367348 9.600019999999985e-05 1.616326530612245 9.699999999999985e-05 1.616326530612245 9.700019999999985e-05 1.683673469387755 9.799999999999985e-05 1.683673469387755 9.800019999999985e-05 1.7510204081632654 9.899999999999984e-05 1.7510204081632654 9.900019999999985e-05 1.8183673469387756 9.999999999999984e-05 1.8183673469387756 0.00010000019999999984 1.8857142857142857 0.00010099999999999984 1.8857142857142857 0.00010100019999999984 1.953061224489796 0.00010199999999999984 1.953061224489796 0.00010200019999999984 2.0204081632653064 0.00010299999999999983 2.0204081632653064 0.00010300019999999983 2.0877551020408163 0.00010399999999999983 2.0877551020408163 0.00010400019999999983 2.1551020408163266 0.00010499999999999983 2.1551020408163266 0.00010500019999999983 2.222448979591837 0.00010599999999999983 2.222448979591837 0.00010600019999999983 2.289795918367347 0.00010699999999999982 2.289795918367347 0.00010700019999999982 2.357142857142857 0.00010799999999999982 2.357142857142857 0.00010800019999999982 2.4244897959183676 0.00010899999999999982 2.4244897959183676 0.00010900019999999982 2.4918367346938775 0.00010999999999999981 2.4918367346938775 0.00011000019999999981 2.559183673469388 0.00011099999999999981 2.559183673469388 0.00011100019999999981 2.626530612244898 0.00011199999999999981 2.626530612244898 0.00011200019999999981 2.6938775510204085 0.0001129999999999998 2.6938775510204085 0.0001130001999999998 2.7612244897959184 0.0001139999999999998 2.7612244897959184 0.0001140001999999998 2.8285714285714287 0.0001149999999999998 2.8285714285714287 0.0001150001999999998 2.895918367346939 0.0001159999999999998 2.895918367346939 0.0001160001999999998 2.963265306122449 0.0001169999999999998 2.963265306122449 0.0001170001999999998 3.0306122448979593 0.00011799999999999979 3.0306122448979593 0.00011800019999999979 3.0979591836734697 0.00011899999999999979 3.0979591836734697 0.00011900019999999979 3.1653061224489796 0.00011999999999999979 3.1653061224489796 0.00012000019999999979 3.23265306122449 0.00012099999999999978 3.23265306122449 0.00012100019999999978 3.3 0.00012199999999999978 3.3)
V12 __VREG_s 0 DC 1 PWL(0 1 1.1e-05 1 1.10002e-05 1 1.2e-05 1 1.20002e-05 1 1.3000000000000001e-05 1 1.3000200000000001e-05 1 1.4000000000000001e-05 1 1.4000200000000002e-05 1 1.5000000000000002e-05 1 1.5000200000000003e-05 1 1.6000000000000003e-05 1 1.6000200000000003e-05 1 1.7000000000000003e-05 1 1.7000200000000004e-05 1 1.8000000000000004e-05 1 1.8000200000000004e-05 1 1.9000000000000004e-05 1 1.9000200000000005e-05 1 2.0000000000000005e-05 1 2.0000200000000005e-05 1 2.1000000000000006e-05 1 2.1000200000000006e-05 1 2.2000000000000006e-05 1 2.2000200000000007e-05 1 2.3000000000000007e-05 1 2.3000200000000007e-05 1 2.4000000000000007e-05 1 2.4000200000000008e-05 1 2.5000000000000008e-05 1 2.500020000000001e-05 1 2.600000000000001e-05 1 2.600020000000001e-05 1 2.700000000000001e-05 1 2.700020000000001e-05 1 2.800000000000001e-05 1 2.800020000000001e-05 1 2.900000000000001e-05 1 2.900020000000001e-05 1 3.000000000000001e-05 1 3.000020000000001e-05 1 3.100000000000001e-05 1 3.100020000000001e-05 1 3.2000000000000005e-05 1 3.2000200000000006e-05 1 3.3e-05 1 3.30002e-05 1 3.4e-05 1 3.40002e-05 1 3.5e-05 1 3.50002e-05 1 3.5999999999999994e-05 1 3.6000199999999995e-05 1 3.699999999999999e-05 1 3.700019999999999e-05 1 3.799999999999999e-05 1 3.800019999999999e-05 1 3.8999999999999986e-05 1 3.9000199999999986e-05 1 3.999999999999998e-05 1 4.000019999999998e-05 1 4.099999999999998e-05 1 4.100019999999998e-05 1 4.199999999999998e-05 1 4.200019999999998e-05 1 4.2999999999999975e-05 1 4.3000199999999975e-05 1 4.399999999999997e-05 1 4.400019999999997e-05 1 4.499999999999997e-05 1 4.500019999999997e-05 1 4.5999999999999966e-05 1 4.6000199999999967e-05 1 4.699999999999996e-05 1 4.7000199999999964e-05 1 4.799999999999996e-05 1 4.800019999999996e-05 1 4.899999999999996e-05 1 4.900019999999996e-05 1 4.9999999999999955e-05 1 5.0000199999999955e-05 1 5.099999999999995e-05 1 5.100019999999995e-05 1 5.199999999999995e-05 1 5.200019999999995e-05 1 5.2999999999999947e-05 1 5.300019999999995e-05 1 5.3999999999999944e-05 1 5.4000199999999944e-05 1 5.499999999999994e-05 1 5.500019999999994e-05 1 5.599999999999994e-05 1 5.600019999999994e-05 1 5.6999999999999935e-05 1 5.7000199999999936e-05 1 5.799999999999993e-05 1 5.800019999999993e-05 1 5.899999999999993e-05 1 5.900019999999993e-05 1 5.999999999999993e-05 1 6.000019999999993e-05 1 6.0999999999999924e-05 1 6.1000199999999925e-05 1 7.199999999999992e-05 1 7.200019999999992e-05 1 7.299999999999992e-05 1 7.300019999999992e-05 1 7.399999999999991e-05 1 7.400019999999992e-05 1 7.499999999999991e-05 1 7.500019999999991e-05 1 7.599999999999991e-05 1 7.600019999999991e-05 1 7.69999999999999e-05 1 7.700019999999991e-05 1 7.79999999999999e-05 1 7.80001999999999e-05 1 7.89999999999999e-05 1 7.90001999999999e-05 1 7.99999999999999e-05 1 8.00001999999999e-05 1 8.09999999999999e-05 1 8.10001999999999e-05 1 8.199999999999989e-05 1 8.200019999999989e-05 1 8.299999999999989e-05 1 8.300019999999989e-05 1 8.399999999999989e-05 1 8.400019999999989e-05 1 8.499999999999988e-05 1 8.500019999999988e-05 1 8.599999999999988e-05 1 8.600019999999988e-05 1 8.699999999999988e-05 1 8.700019999999988e-05 1 8.799999999999988e-05 1 8.800019999999988e-05 1 8.899999999999987e-05 1 8.900019999999987e-05 1 8.999999999999987e-05 1 9.000019999999987e-05 1 9.099999999999987e-05 1 9.100019999999987e-05 1 9.199999999999986e-05 1 9.200019999999986e-05 1 9.299999999999986e-05 1 9.300019999999986e-05 1 9.399999999999986e-05 1 9.400019999999986e-05 1 9.499999999999986e-05 1 9.500019999999986e-05 1 9.599999999999985e-05 1 9.600019999999985e-05 1 9.699999999999985e-05 1 9.700019999999985e-05 1 9.799999999999985e-05 1 9.800019999999985e-05 1 9.899999999999984e-05 1 9.900019999999985e-05 1 9.999999999999984e-05 1 0.00010000019999999984 1 0.00010099999999999984 1 0.00010100019999999984 1 0.00010199999999999984 1 0.00010200019999999984 1 0.00010299999999999983 1 0.00010300019999999983 1 0.00010399999999999983 1 0.00010400019999999983 1 0.00010499999999999983 1 0.00010500019999999983 1 0.00010599999999999983 1 0.00010600019999999983 1 0.00010699999999999982 1 0.00010700019999999982 1 0.00010799999999999982 1 0.00010800019999999982 1 0.00010899999999999982 1 0.00010900019999999982 1 0.00010999999999999981 1 0.00011000019999999981 1 0.00011099999999999981 1 0.00011100019999999981 1 0.00011199999999999981 1 0.00011200019999999981 1 0.0001129999999999998 1 0.0001130001999999998 1 0.0001139999999999998 1 0.0001140001999999998 1 0.0001149999999999998 1 0.0001150001999999998 1 0.0001159999999999998 1 0.0001160001999999998 1 0.0001169999999999998 1 0.0001170001999999998 1 0.00011799999999999979 1 0.00011800019999999979 1 0.00011899999999999979 1 0.00011900019999999979 1 0.00011999999999999979 1 0.00012000019999999979 1 0.00012099999999999978 1 0.00012100019999999978 1 0.00012199999999999978 1)
X13 __VREF_v VREF __VREF_s 0 inout_sw_mod
V14 __VREF_v 0 DC 1.6 PWL(0 1.6 9.999999999999999e-06 1.6 1.00002e-05 1.6 6.0999999999999924e-05 1.6 6.1000199999999925e-05 1.6 7.099999999999992e-05 1.6 7.100019999999992e-05 1.6 0.00012199999999999978 1.6)
V15 __VREF_s 0 DC 1 PWL(0 1 9.999999999999999e-06 1 1.00002e-05 1 6.0999999999999924e-05 1 6.1000199999999925e-05 1 7.099999999999992e-05 1 7.100019999999992e-05 1 0.00012199999999999978 1)
.tran 10e-9 0.00012199999999999978
.control
run
set filetype=binary
write
exit
.endc
.probe V(outn) V(VREG) V(vgnd) V(vpwr) V(VREF) V(CLK) V(outp)
.end
